`define D_INIT_FILE "dmem.hex"
`define I_INIT_FILE "imem.hex"
