`define D_INIT_FILE "/home/yc/proj/1_TFLM/sw/build/dmem.hex"
`define I_INIT_FILE "/home/yc/proj/1_TFLM/sw/build/imem.hex"
